module main

fn internal_word_list() []string {
	return [
		'the',
		'for',
		'use',
		'anyone',
		'anywhere',
		'cost',
		'and',
		'with',
		'almost',
		'whatsoever',
		'may',
		'copy',
		'give',
		'away',
		'under',
		'terms',
		'included',
		'this',
		'online',
		'updated',
		'set',
		'encoding',
		'cover',
		'took',
		'his',
		'bottle',
		'from',
		'corner',
		'hypodermic',
		'syringe',
		'its',
		'neat',
		'morocco',
		'case',
		'long',
		'white',
		'nervous',
		'fingers',
		'adjusted',
		'delicate',
		'needle',
		'rolled',
		'back',
		'left',
		'some',
		'little',
		'time',
		'eyes',
		'rested',
		'upon',
		'sinewy',
		'forearm',
		'wrist',
		'all',
		'dotted',
		'scarred',
		'thrust',
		'sharp',
		'point',
		'home',
		'pressed',
		'down',
		'tiny',
		'piston',
		'sank',
		'into',
		'sigh',
		'times',
		'day',
		'many',
		'months',
		'had',
		'witnessed',
		'but',
		'custom',
		'not',
		'reconciled',
		'mind',
		'contrary',
		'become',
		'more',
		'irritable',
		'sight',
		'conscience',
		'swelled',
		'nightly',
		'within',
		'thought',
		'that',
		'lacked',
		'courage',
		'protest',
		'again',
		'registered',
		'vow',
		'should',
		'deliver',
		'soul',
		'subject',
		'there',
		'was',
		'cool',
		'nonchalant',
		'air',
		'companion',
		'which',
		'made',
		'him',
		'last',
		'man',
		'whom',
		'one',
		'would',
		'care',
		'take',
		'anything',
		'liberty',
		'great',
		'powers',
		'masterly',
		'manner',
		'experience',
		'qualities',
		'diffident',
		'backward',
		'crossing',
		'afternoon',
		'whether',
		'taken',
		'lunch',
		'additional',
		'produced',
		'extreme',
		'suddenly',
		'felt',
		'could',
		'hold',
		'out',
		'longer',
		'raised',
		'languidly',
		'old',
		'volume',
		'opened',
		'cocaine',
		'solution',
		'you',
		'try',
		'indeed',
		'answered',
		'brusquely',
		'has',
		'got',
		'over',
		'campaign',
		'yet',
		'cannot',
		'afford',
		'throw',
		'any',
		'extra',
		'strain',
		'smiled',
		'vehemence',
		'are',
		'right',
		'said',
		'suppose',
		'influence',
		'physically',
		'bad',
		'find',
		'however',
		'clarifying',
		'secondary',
		'action',
		'matter',
		'small',
		'moment',
		'earnestly',
		'brain',
		'say',
		'roused',
		'excited',
		'morbid',
		'process',
		'involves',
		'increased',
		'leave',
		'permanent',
		'weakness',
		'know',
		'too',
		'what',
		'black',
		'reaction',
		'comes',
		'game',
		'hardly',
		'worth',
		'candle',
		'mere',
		'passing',
		'pleasure',
		'risk',
		'loss',
		'those',
		'have',
		'been',
		'speak',
		'only',
		'comrade',
		'another',
		'medical',
		'whose',
		'extent',
		'answerable',
		'did',
		'seem',
		'offended',
		'put',
		'together',
		'leaned',
		'elbows',
		'arms',
		'chair',
		'like',
		'who',
		'relish',
		'rebels',
		'stagnation',
		'problems',
		'work',
		'most',
		'abstruse',
		'cryptogram',
		'intricate',
		'analysis',
		'own',
		'proper',
		'atmosphere',
		'can',
		'dispense',
		'then',
		'artificial',
		'stimulants',
		'abhor',
		'dull',
		'routine',
		'existence',
		'crave',
		'mental',
		'exaltation',
		'why',
		'chosen',
		'particular',
		'rather',
		'created',
		'world',
		'unofficial',
		'raising',
		'eyebrows',
		'consulting',
		'detective',
		'highest',
		'court',
		'appeal',
		'detection',
		'their',
		'way',
		'normal',
		'laid',
		'before',
		'examine',
		'data',
		'expert',
		'pronounce',
		'opinion',
		'claim',
		'credit',
		'such',
		'cases',
		'name',
		'figures',
		'newspaper',
		'itself',
		'finding',
		'field',
		'peculiar',
		'reward',
		'yourself',
		'methods',
		'cordially',
		'never',
		'struck',
		'life',
		'even',
		'embodied',
		'brochure',
		'somewhat',
		'fantastic',
		'title',
		'shook',
		'head',
		'sadly',
		'glanced',
		'ought',
		'exact',
		'science',
		'treated',
		'same',
		'cold',
		'attempted',
		'tinge',
		'produces',
		'much',
		'effect',
		'worked',
		'elopement',
		'fifth',
		'romance',
		'tamper',
		'facts',
		'suppressed',
		'least',
		'just',
		'sense',
		'proportion',
		'observed',
		'treating',
		'them',
		'deserved',
		'mention',
		'curious',
		'analytical',
		'reasoning',
		'effects',
		'causes',
		'succeeded',
		'unraveling',
		'annoyed',
		'criticism',
		'specially',
		'designed',
		'please',
		'confess',
		'irritated',
		'egotism',
		'seemed',
		'demand',
		'every',
		'line',
		'pamphlet',
		'devoted',
		'special',
		'doings',
		'than',
		'once',
		'during',
		'years',
		'lived',
		'vanity',
		'underlay',
		'quiet',
		'didactic',
		'remark',
		'sat',
		'nursing',
		'wounded',
		'leg',
		'bullet',
		'through',
		'though',
		'prevent',
		'walking',
		'ached',
		'wearily',
		'change',
		'weather',
		'practice',
		'extended',
		'recently',
		'after',
		'while',
		'filling',
		'pipe',
		'consulted',
		'week',
		'probably',
		'come',
		'front',
		'lately',
		'service',
		'power',
		'quick',
		'intuition',
		'deficient',
		'wide',
		'range',
		'knowledge',
		'essential',
		'higher',
		'art',
		'concerned',
		'will',
		'possessed',
		'features',
		'interest',
		'able',
		'refer',
		'two',
		'parallel',
		'other',
		'suggested',
		'true',
		'letter',
		'morning',
		'assistance',
		'tossed',
		'spoke',
		'crumpled',
		'sheet',
		'foreign',
		'notepaper',
		'catching',
		'profusion',
		'notes',
		'admiration',
		'stray',
		'testifying',
		'ardent',
		'speaks',
		'pupil',
		'master',
		'rates',
		'highly',
		'lightly',
		'gifts',
		'himself',
		'possesses',
		'three',
		'necessary',
		'ideal',
		'deduction',
		'wanting',
		'now',
		'works',
		'cried',
		'laughing',
		'guilty',
		'several',
		'monographs',
		'technical',
		'subjects',
		'example',
		'between',
		'enumerate',
		'hundred',
		'forty',
		'forms',
		'coloured',
		'plates',
		'difference',
		'ash',
		'turning',
		'criminal',
		'trials',
		'sometimes',
		'supreme',
		'importance',
		'clue',
		'definitely',
		'murder',
		'done',
		'smoking',
		'lunkah',
		'obviously',
		'narrows',
		'your',
		'search',
		'trained',
		'eye',
		'fluff',
		'cabbage',
		'potato',
		'genius',
		'remarked',
		'appreciate',
		'monograph',
		'tracing',
		'footsteps',
		'remarks',
		'uses',
		'plaster',
		'preserver',
		'impresses',
		'trade',
		'form',
		'hand',
		'lithotypes',
		'hands',
		'slaters',
		'sailors',
		'weavers',
		'practical',
		'scientific',
		'unclaimed',
		'bodies',
		'criminals',
		'weary',
		'hobby',
		'greatest',
		'especially',
		'since',
		'observing',
		'implies',
		'leaning',
		'sending',
		'thick',
		'blue',
		'wreaths',
		'shows',
		'lets',
		'when',
		'dispatched',
		'telegram',
		'both',
		'see',
		'how',
		'arrived',
		'sudden',
		'impulse',
		'part',
		'mentioned',
		'simplicity',
		'chuckling',
		'absurdly',
		'simple',
		'serve',
		'define',
		'limits',
		'tells',
		'reddish',
		'mould',
		'adhering',
		'instep',
		'opposite',
		'they',
		'pavement',
		'thrown',
		'earth',
		'lies',
		'difficult',
		'avoid',
		'treading',
		'entering',
		'tint',
		'found',
		'far',
		'nowhere',
		'else',
		'rest',
		'deduce',
		'course',
		'knew',
		'written',
		'also',
		'open',
		'desk',
		'stamps',
		'bundle',
		'send',
		'factors',
		'remains',
		'must',
		'truth',
		'certainly',
		'replied',
		'thing',
		'simplest',
		'think',
		'were',
		'theories',
		'severe',
		'taking',
		'second',
		'dose',
		'delighted',
		'look',
		'problem',
		'might',
		'submit',
		'heard',
		'object',
		'daily',
		'without',
		'leaving',
		'impress',
		'observer',
		'read',
		'here',
		'watch',
		'possession',
		'kindness',
		'let',
		'character',
		'habits',
		'late',
		'handed',
		'slight',
		'feeling',
		'amusement',
		'heart',
		'test',
		'impossible',
		'intended',
		'lesson',
		'against',
		'dogmatic',
		'tone',
		'assumed',
		'balanced',
		'gazed',
		'hard',
		'dial',
		'examined',
		'first',
		'naked',
		'powerful',
		'convex',
		'lens',
		'keep',
		'smiling',
		'face',
		'finally',
		'snapped',
		'cleaned',
		'robs',
		'suggestive',
		'being',
		'sent',
		'accused',
		'putting',
		'forward',
		'lame',
		'impotent',
		'excuse',
		'failure',
		'expect',
		'uncleaned',
		'research',
		'entirely',
		'barren',
		'staring',
		'ceiling',
		'dreamy',
		'correction',
		'judge',
		'belonged',
		'elder',
		'brother',
		'inherited',
		'father',
		'gather',
		'doubt',
		'suggests',
		'date',
		'nearly',
		'fifty',
		'initials',
		'generation',
		'usually',
		'descends',
		'eldest',
		'son',
		'likely',
		'remember',
		'dead',
		'therefore',
		'untidy',
		'careless',
		'good',
		'prospects',
		'threw',
		'chances',
		'poverty',
		'occasional',
		'short',
		'intervals',
		'prosperity',
		'drink',
		'died',
		'sprang',
		'limped',
		'about',
		'room',
		'bitterness',
		'unworthy',
		'believed',
		'descended',
		'inquires',
		'history',
		'unhappy',
		'pretend',
		'fanciful',
		'believe',
		'unkind',
		'plainly',
		'touch',
		'dear',
		'doctor',
		'kindly',
		'pray',
		'accept',
		'apologies',
		'abstract',
		'forgotten',
		'personal',
		'painful',
		'assure',
		'until',
		'wonderful',
		'get',
		'these',
		'absolutely',
		'correct',
		'luck',
		'balance',
		'accurate',
		'guess',
		'shocking',
		'logical',
		'faculty',
		'seems',
		'strange',
		'because',
		'follow',
		'train',
		'observe',
		'large',
		'inferences',
		'depend',
		'began',
		'stating',
		'lower',
		'notice',
		'dinted',
		'places',
		'cut',
		'marked',
		'habit',
		'keeping',
		'objects',
		'coins',
		'keys',
		'pocket',
		'feat',
		'assume',
		'treats',
		'cavalierly',
		'very',
		'inference',
		'inherits',
		'article',
		'value',
		'pretty',
		'well',
		'provided',
		'respects',
		'nodded',
		'show',
		'followed',
		'customary',
		'scratch',
		'number',
		'ticket',
		'inside',
		'handy',
		'label',
		'lost',
		'transposed',
		'less',
		'four',
		'numbers',
		'visible',
		'often',
		'low',
		'water',
		'bursts',
		'redeemed',
		'pledge',
		'ask',
		'inner',
		'plate',
		'contains',
		'thousands',
		'scratches',
		'round',
		'where',
		'key',
		'slipped',
		'sober',
		'scored',
		'winds',
		'night',
		'leaves',
		'traces',
		'unsteady',
		'mystery',
		'clear',
		'daylight',
		'regret',
		'injustice',
		'faith',
		'marvellous',
		'inquiry',
		'foot',
		'live',
		'window',
		'ever',
		'dreary',
		'dismal',
		'yellow',
		'fog',
		'swirls',
		'street',
		'drifts',
		'across',
		'houses',
		'hopelessly',
		'prosaic',
		'having',
		'exert',
		'save',
		'function',
		'mouth',
		'reply',
		'tirade',
		'crisp',
		'knock',
		'our',
		'landlady',
		'entered',
		'bearing',
		'card',
		'brass',
		'salver',
		'young',
		'lady',
		'sir',
		'she',
		'addressing',
		'step',
		'prefer',
		'remain',
		'firm',
		'outward',
		'composure',
		'blonde',
		'dainty',
		'gloved',
		'dressed',
		'perfect',
		'taste',
		'plainness',
		'her',
		'costume',
		'bore',
		'suggestion',
		'limited',
		'means',
		'dress',
		'sombre',
		'greyish',
		'beige',
		'untrimmed',
		'unbraided',
		'wore',
		'turban',
		'hue',
		'relieved',
		'suspicion',
		'feather',
		'side',
		'neither',
		'regularity',
		'feature',
		'nor',
		'beauty',
		'complexion',
		'expression',
		'sweet',
		'amiable',
		'singularly',
		'spiritual',
		'women',
		'extends',
		'nations',
		'separate',
		'continents',
		'looked',
		'gave',
		'clearer',
		'promise',
		'refined',
		'sensitive',
		'nature',
		'seat',
		'placed',
		'lip',
		'trembled',
		'quivered',
		'showed',
		'sign',
		'intense',
		'inward',
		'agitation',
		'enabled',
		'employer',
		'unravel',
		'domestic',
		'impressed',
		'skill',
		'repeated',
		'mine',
		'imagine',
		'utterly',
		'situation',
		'myself',
		'rubbed',
		'glistened',
		'hawklike',
		'brisk',
		'business',
		'tones',
		'position',
		'sure',
		'rising',
		'surprise',
		'held',
		'detain',
		'friend',
		'enough',
		'stop',
		'relapsed',
		'continued',
		'officer',
		'regiment',
		'quite',
		'child',
		'mother',
		'relative',
		'boarding',
		'remained',
		'seventeen',
		'age',
		'year',
		'senior',
		'captain',
		'obtained',
		'twelve',
		'came',
		'safe',
		'directed',
		'giving',
		'address',
		'message',
		'full',
		'love',
		'reaching',
		'drove',
		'informed',
		'staying',
		'gone',
		'returned',
		'waited',
		'news',
		'advice',
		'manager',
		'hotel',
		'police',
		'next',
		'advertised',
		'papers',
		'inquiries',
		'led',
		'word',
		'hope',
		'peace',
		'comfort',
		'throat',
		'choking',
		'sob',
		'sentence',
		'asked',
		'opening',
		'ten',
		'ago',
		'nothing',
		'suggest',
		'clothes',
		'books',
		'officers',
		'charge',
		'friends',
		'major',
		'retired',
		'singular',
		'described',
		'six',
		'appeared',
		'asking',
		'advantage',
		'appended',
		'family',
		'capacity',
		'governess',
		'published',
		'column',
		'post',
		'box',
		'addressed',
		'contain',
		'lustrous',
		'pearl',
		'writing',
		'enclosed',
		'always',
		'similar',
		'containing',
		'sender',
		'pronounced',
		'rare',
		'variety',
		'yourselves',
		'handsome',
		'flat',
		'finest',
		'pearls',
		'seen',
		'statement',
		'occurred',
		'later',
		'received',
		'perhaps',
		'envelope',
		'postman',
		'quality',
		'paper',
		'sixpence',
		'packet',
		'stationery',
		'third',
		'pillar',
		'outside',
		'seven',
		'bring',
		'wronged',
		'woman',
		'shall',
		'justice',
		'vain',
		'unknown',
		'really',
		'intend',
		'exactly',
		'want',
		'says',
		'something',
		'appealing',
		'voice',
		'proud',
		'happy',
		'fervently',
		'kind',
		'producing',
		'half',
		'dozen',
		'pieces',
		'model',
		'client',
		'spread',
		'table',
		'darting',
		'glances',
		'disguised',
		'except',
		'presently',
		'question',
		'authorship',
		'break',
		'twirl',
		'final',
		'person',
		'false',
		'hopes',
		'unlike',
		'expected',
		'hear',
		'allow',
		'visitor',
		'bright',
		'glance',
		'replaced',
		'bosom',
		'hurried',
		'watched',
		'briskly',
		'grey',
		'speck',
		'crowd',
		'attractive',
		'exclaimed',
		'lit',
		'drooping',
		'eyelids',
		'positively',
		'inhuman',
		'gently',
		'judgment',
		'biased',
		'factor',
		'emotional',
		'winning',
		'hanged',
		'poisoning',
		'children',
		'repellant',
		'spent',
		'quarter',
		'million',
		'poor',
		'make',
		'exceptions',
		'exception',
		'disproves',
		'rule',
		'occasion',
		'study',
		'legible',
		'regular',
		'force',
		'letters',
		'rise',
		'above',
		'common',
		'herd',
		'illegibly',
		'write',
		'capitals',
		'going',
		'few',
		'references',
		'recommend',
		'remarkable',
		'penned',
		'hour',
		'thoughts',
		'daring',
		'writer',
		'ran',
		'smiles',
		'deep',
		'rich',
		'overhung',
		'youth',
		'sobered',
		'mused',
		'dangerous',
		'plunged',
		'furiously',
		'latest',
		'treatise',
		'pathology',
		'army',
		'surgeon',
		'weak',
		'weaker',
		'dare',
		'unit',
		'future',
		'better',
		'surely',
		'attempt',
		'brighten',
		'five',
		'eager',
		'excellent',
		'mood',
		'alternated',
		'fits',
		'blackest',
		'depression',
		'cup',
		'tea',
		'poured',
		'appear',
		'admit',
		'solved',
		'discovered',
		'fact',
		'details',
		'still',
		'added',
		'files',
		'obtuse',
		'fail',
		'disappears',
		'visited',
		'denies',
		'dies',
		'daughter',
		'receives',
		'valuable',
		'present',
		'culminates',
		'describes',
		'wrong',
		'presents',
		'begin',
		'death',
		'unless',
		'heir',
		'knows',
		'desires',
		'theory',
		'meet',
		'strangely',
		'alive',
		'pensively',
		'expedition',
		'solve',
		'past',
		'picked',
		'hat',
		'heaviest',
		'stick',
		'revolver',
		'drawer',
		'serious',
		'muffled',
		'dark',
		'cloak',
		'composed',
		'pale',
		'feel',
		'uneasiness',
		'enterprise',
		'embarking',
		'readily',
		'questions',
		'allusions',
		'papa',
		'command',
		'troops',
		'deal',
		'understand',
		'slightest',
		'brought',
		'unfolded',
		'carefully',
		'smoothed',
		'knee',
		'double',
		'native',
		'pinned',
		'board',
		'diagram',
		'appears',
		'plan',
		'building',
		'numerous',
		'halls',
		'corridors',
		'passages',
		'cross',
		'red',
		'ink',
		'faded',
		'crosses',
		'touching',
		'rough',
		'coarse',
		'characters',
		'bears',
		'evidently',
		'document',
		'kept',
		'clean',
		'prove',
		'suspect',
		'turn',
		'deeper',
		'subtle',
		'supposed',
		'reconsider',
		'ideas',
		'cab',
		'drawn',
		'brow',
		'vacant',
		'thinking',
		'intently',
		'chatted',
		'undertone',
		'possible',
		'outcome',
		'maintained',
		'reserve',
		'end',
		'journey',
		'evening',
		'dense',
		'drizzly',
		'lay',
		'city',
		'clouds',
		'drooped',
		'muddy',
		'streets',
		'lamps',
		'misty',
		'splotches',
		'diffused',
		'light',
		'feeble',
		'circular',
		'glimmer',
		'slimy',
		'glare',
		'streamed',
		'steamy',
		'vaporous',
		'murky',
		'shifting',
		'radiance',
		'crowded',
		'eerie',
		'endless',
		'procession',
		'faces',
		'flitted',
		'narrow',
		'bars',
		'glad',
		'haggard',
		'merry',
		'human',
		'gloom',
		'heavy',
		'engaged',
		'combined',
		'depressed',
		'suffering',
		'alone',
		'superior',
		'petty',
		'influences',
		'jotted',
		'memoranda',
		'crowds',
		'already',
		'continuous',
		'stream',
		'hansoms',
		'rattling',
		'cargoes',
		'men',
		'beshawled',
		'reached',
		'rendezvous',
		'coachman',
		'accosted',
		'parties',
		'gentlemen',
		'bent',
		'pair',
		'miss',
		'certain',
		'dogged',
		'companions',
		'shrill',
		'whistle',
		'door',
		'mounted',
		'driver',
		'whipped',
		'horse',
		'furious',
		'pace',
		'foggy',
		'driving',
		'place',
		'errand',
		'invitation',
		'either',
		'complete',
		'reason',
		'important',
		'issues',
		'hang',
		'demeanor',
		'resolute',
		'collected',
		'endeavored',
		'cheer',
		'amuse',
		'adventures',
		'tell',
		'stories',
		'slightly',
		'involved',
		'declares',
		'told',
		'moving',
		'anecdote',
		'musket',
		'tent',
		'fired',
		'tiger',
		'cub',
		'idea',
		'direction',
		'soon',
		'bearings',
		'fault',
		'muttered',
		'names',
		'rattled',
		'squares',
		'tortuous',
		'making',
		'apparently',
		'bridge',
		'catch',
		'glimpses',
		'river',
		'fleeting',
		'view',
		'stretch',
		'shining',
		'broad',
		'silent',
		'dashed',
		'labyrinth',
		'quest',
		'does',
		'regions',
		'forbidding',
		'lines',
		'brick',
		'tawdry',
		'brilliancy',
		'public',
		'rows',
		'villas',
		'each',
		'fronting',
		'miniature',
		'garden',
		'new',
		'monster',
		'tentacles',
		'giant',
		'throwing',
		'country',
		'drew',
		'house',
		'terrace',
		'inhabited',
		'stopped',
		'neighbours',
		'single',
		'kitchen',
		'knocking',
		'instantly',
		'servant',
		'clad',
		'sash',
		'figure',
		'framed',
		'doorway',
		'suburban',
		'awaits',
		'high',
		'piping',
		'khitmutgar',
		'straight',
		'sordid',
		'passage',
		'worse',
		'furnished',
		'blaze',
		'centre',
		'stood',
		'bristle',
		'hair',
		'fringe',
		'bald',
		'scalp',
		'shot',
		'among',
		'writhed',
		'perpetual',
		'jerk',
		'scowling',
		'instant',
		'repose',
		'given',
		'pendulous',
		'irregular',
		'teeth',
		'strove',
		'feebly',
		'conceal',
		'constantly',
		'spite',
		'obtrusive',
		'baldness',
		'impression',
		'turned',
		'thirtieth',
		'repeating',
		'thin',
		'sanctum',
		'liking',
		'oasis',
		'howling',
		'desert',
		'astonished',
		'appearance',
		'apartment',
		'invited',
		'sorry',
		'diamond',
		'setting',
		'richest',
		'glossiest',
		'curtains',
		'tapestries',
		'draped',
		'walls',
		'looped',
		'expose',
		'painting',
		'vase',
		'carpet',
		'soft',
		'pleasantly',
		'bed',
		'moss',
		'athwart',
		'luxury',
		'huge',
		'hookah',
		'mat',
		'lamp',
		'fashion',
		'silver',
		'dove',
		'hung',
		'invisible',
		'golden',
		'wire',
		'burned',
		'filled',
		'aromatic',
		'odour',
		'jerking',
		'grave',
		'doubts',
		'mitral',
		'valve',
		'aortic',
		'rely',
		'listened',
		'requested',
		'unable',
		'amiss',
		'ecstasy',
		'fear',
		'shivered',
		'cause',
		'anxiety',
		'airily',
		'sufferer',
		'suspicions',
		'refrained',
		'hot',
		'callous',
		'reference',
		'grew',
		'lips',
		'whatever',
		'escort',
		'witnesses',
		'bold',
		'officials',
		'settle',
		'everything',
		'ourselves',
		'annoy',
		'publicity',
		'settee',
		'blinked',
		'watery',
		'choose',
		'further',
		'agreement',
		'offer',
		'glass',
		'wines',
		'trust',
		'objection',
		'mild',
		'balsamic',
		'tobacco',
		'invaluable',
		'sedative',
		'applied',
		'taper',
		'bowl',
		'smoke',
		'bubbled',
		'merrily',
		'heads',
		'advanced',
		'chins',
		'jerky',
		'fellow',
		'puffed',
		'uneasily',
		'determined',
		'feared',
		'disregard',
		'request',
		'unpleasant',
		'people',
		'confidence',
		'discretion',
		'orders',
		'proceed',
		'retiring',
		'tastes',
		'policeman',
		'natural',
		'shrinking',
		'seldom',
		'contact',
		'elegance',
		'around',
		'call',
		'patron',
		'arts',
		'landscape',
		'genuine',
		'partial',
		'modern',
		'school',
		'learn',
		'desire',
		'interview',
		'best',
		'angry',
		'words',
		'terrible',
		'start',
		'ventured',
		'laughed',
		'ears',
		'prepare',
		'showing',
		'stand',
		'points',
		'story',
		'ignorant',
		'guessed',
		'eleven',
		'prospered',
		'sum',
		'money',
		'collection',
		'staff',
		'servants',
		'advantages',
		'bought',
		'sensation',
		'caused',
		'knowing',
		'discussed',
		'freely',
		'presence',
		'used',
		'join',
		'happened',
		'whole',
		'secret',
		'hidden',
		'fate',
		'positive',
		'fearful',
		'employed',
		'act',
		'porters',
		'champion',
		'aversion',
		'wooden',
		'legs',
		'actually',
		'proved',
		'harmless',
		'tradesman',
		'canvassing',
		'pay',
		'hush',
		'whim',
		'events',
		'shock',
		'fainted',
		'sickened',
		'discover',
		'scrawling',
		'suffered',
		'enlarged',
		'spleen',
		'became',
		'rapidly',
		'towards',
		'beyond',
		'wished',
		'propped',
		'pillows',
		'breathing',
		'heavily',
		'besought',
		'lock',
		'grasping',
		'broken',
		'emotion',
		'pain',
		'weighs',
		'treatment',
		'orphan',
		'cursed',
		'greed',
		'besetting',
		'sin',
		'withheld',
		'treasure',
		'hers',
		'blind',
		'foolish',
		'avarice',
		'bear',
		'share',
		'chaplet',
		'dipped',
		'beside',
		'although',
		'design',
		'sons',
		'fair',
		'recovered',
		'concealed',
		'chain',
		'arrival',
		'walked',
		'station',
		'admitted',
		'faithful',
		'division',
		'heated',
		'sprung',
		'paroxysm',
		'anger',
		'dusky',
		'fell',
		'backwards',
		'cutting',
		'stooped',
		'horror',
		'distracted',
		'wondering',
		'recognise',
		'chance',
		'quarrel',
		'gash',
		'official',
		'bringing',
		'anxious',
		'necessity',
		'pondering',
		'looking',
		'saw',
		'stole',
		'bolted',
		'behind',
		'need',
		'killed',
		'hide',
		'kill',
		'blow',
		'sealed',
		'asleep',
		'decide',
		'innocence',
		'tradesmen',
		'disposed',
		'body',
		'days',
		'mysterious',
		'blamed',
		'clung',
		'wish',
		'horrible',
		'stared',
		'wildly',
		'jaw',
		'dropped',
		'yelled',
		'forget',
		'sake',
		'gaze',
		'fixed',
		'darkness',
		'whitening',
		'nose',
		'bearded',
		'hairy',
		'wild',
		'cruel',
		'rushed',
		'pulse',
		'ceased',
		'beat',
		'searched',
		'intruder',
		'footmark',
		'trace',
		'conjured',
		'fierce',
		'striking',
		'proof',
		'agencies',
		'cupboards',
		'boxes',
		'rifled',
		'chest',
		'torn',
		'piece',
		'scrawled',
		'phrase',
		'meant',
		'none',
		'property',
		'stolen',
		'naturally',
		'associated',
		'incident',
		'haunted',
		'relight',
		'moments',
		'absorbed',
		'listening',
		'narrative',
		'account',
		'deadly',
		'faint',
		'rallied',
		'drinking',
		'quietly',
		'carafe',
		'abstracted',
		'lids',
		'glittering',
		'complained',
		'bitterly',
		'tax',
		'sagacity',
		'utmost',
		'obvious',
		'pride',
		'puffs',
		'overgrown',
		'spoken',
		'weeks',
		'dug',
		'delved',
		'maddening',
		'splendour',
		'missing',
		'riches',
		'discussion',
		'averse',
		'inclined',
		'parted',
		'gossip',
		'trouble',
		'persuade',
		'detached',
		'destitute',
		'extremely',
		'waved',
		'trustees',
		'altogether',
		'plenty',
		'desired',
		'scurvy',
		'mauvais',
		'things',
		'went',
		'rooms',
		'event',
		'drive',
		'explained',
		'views',
		'welcome',
		'visitors',
		'twitching',
		'luxurious',
		'spring',
		'feet',
		'return',
		'delay',
		'coiled',
		'tube',
		'curtain',
		'befrogged',
		'topcoat',
		'collar',
		'cuffs',
		'buttoned',
		'tightly',
		'closeness',
		'finished',
		'attire',
		'cap',
		'hanging',
		'lappets',
		'covered',
		'mobile',
		'peaky',
		'health',
		'fragile',
		'compelled',
		'awaiting',
		'programme',
		'started',
		'off',
		'rapid',
		'talked',
		'rose',
		'rattle',
		'wheels',
		'clever',
		'conclusion',
		'somewhere',
		'indoors',
		'cubic',
		'space',
		'everywhere',
		'inch',
		'height',
		'adding',
		'heights',
		'allowance',
		'borings',
		'total',
		'seventy',
		'top',
		'knocked',
		'hole',
		'garret',
		'known',
		'resting',
		'rafters',
		'lowered',
		'computes',
		'jewels',
		'sterling',
		'gigantic',
		'secure',
		'rights',
		'needy',
		'heiress',
		'loyal',
		'rejoice',
		'ashamed',
		'lead',
		'stammered',
		'halting',
		'downcast',
		'deaf',
		'babble',
		'clearly',
		'confirmed',
		'dreamily',
		'conscious',
		'pouring',
		'forth',
		'trains',
		'symptoms',
		'imploring',
		'quack',
		'nostrums',
		'leather',
		'answers',
		'overheard',
		'caution',
		'danger',
		'drops',
		'castor',
		'oil',
		'strychnine',
		'doses',
		'pulled',
		'stage',
		'damp',
		'fairly',
		'fine',
		'warm',
		'wind',
		'blew',
		'westward',
		'moved',
		'slowly',
		'sky',
		'moon',
		'peeping',
		'rifts',
		'distance',
		'carriage',
		'grounds',
		'girt',
		'stone',
		'wall',
		'topped',
		'formed',
		'entrance',
		'guide',
		'gruff',
		'grumbling',
		'sound',
		'clanking',
		'jarring',
		'swung',
		'lantern',
		'protruded',
		'twinkling',
		'unexpected',
		'obstacle',
		'perplexed',
		'helpless',
		'guarantee',
		'wait',
		'road',
		'porter',
		'inexorably',
		'yours',
		'pays',
		'duty',
		'yes',
		'genially',
		'amateur',
		'fought',
		'rounds',
		'benefit',
		'roared',
		'mistook',
		'instead',
		'stepped',
		'wasted',
		'aimed',
		'joined',
		'fancy',
		'fails',
		'strict',
		'gravel',
		'path',
		'wound',
		'desolate',
		'clump',
		'square',
		'shadow',
		'moonbeam',
		'glimmered',
		'vast',
		'size',
		'deathly',
		'silence',
		'chill',
		'ill',
		'ease',
		'mistake',
		'distinctly',
		'guard',
		'premises',
		'favourite',
		'moonshine',
		'strikes',
		'glint',
		'sits',
		'waiting',
		'minute',
		'coming',
		'alarmed',
		'circles',
		'flickered',
		'wavered',
		'seized',
		'thumping',
		'hearts',
		'straining',
		'sounded',
		'saddest',
		'pitiful',
		'whimpering',
		'frightened',
		'tall',
		'sway',
		'reiterated',
		'rejoicings',
		'closed',
		'monotone',
		'peered',
		'keenly',
		'cumbered',
		'wondrous',
		'affection',
		'passed',
		'sought',
		'marvelled',
		'instinct',
		'protection',
		'surrounded',
		'looks',
		'moles',
		'loose',
		'sort',
		'hill',
		'near',
		'wonder',
		'burst',
		'running',
		'terror',
		'nerves',
		'blubbering',
		'terrified',
		'pleaded',
		'equal',
		'directions',
		'pacing',
		'scared',
		'restless',
		'picking',
		'soothing',
		'bless',
		'calm',
		'hysterical',
		'sorely',
		'tried',
		'patted',
		'murmured',
		'womanly',
		'colour',
		'bloodless',
		'cheeks',
		'locked',
		'answer',
		'likes',
		'peeped',
		'joy',
		'sorrow',
		'chattering',
		'shaken',
		'pass',
		'arm',
		'stairs',
		'knees',
		'trembling',
		'ascended',
		'marks',
		'shapeless',
		'smudges',
		'dust',
		'matting',
		'served',
		'holding',
		'shooting',
		'keen',
		'flight',
		'ended',
		'length',
		'picture',
		'tapestry',
		'doors',
		'along',
		'slow',
		'methodical',
		'close',
		'heels',
		'shadows',
		'streaming',
		'corridor',
		'seeking',
		'receiving',
		'handle',
		'bolt',
		'intaking',
		'breath',
		'devilish',
		'recoiled',
		'vague',
		'shifty',
		'suspended',
		'beneath',
		'smile',
		'unnatural',
		'grin',
		'moonlit',
		'scowl',
		'contortion',
		'recalled',
		'twins',
		'springing',
		'weight',
		'creaked',
		'groaned',
		'yield',
		'flung',
		'snap',
		'chamber',
		'fitted',
		'chemical',
		'laboratory',
		'bottles',
		'littered',
		'burners',
		'retorts',
		'corners',
		'carboys',
		'acid',
		'wicker',
		'baskets',
		'leak',
		'liquid',
		'trickled',
		'peculiarly',
		'pungent',
		'steps',
		'midst',
		'litter',
		'lath',
		'coil',
		'rope',
		'carelessly',
		'seated',
		'heap',
		'sunk',
		'shoulder',
		'ghastly',
		'stiff',
		'hours',
		'limbs',
		'twisted',
		'brown',
		'hammer',
		'rudely',
		'lashed',
		'twine',
		'thrill',
		'stooping',
		'pointed',
		'thorn',
		'stuck',
		'skin',
		'ear',
		'pick',
		'careful',
		'poisoned',
		'finger',
		'thumb',
		'mark',
		'blood',
		'puncture',
		'insoluble',
		'grows',
		'darker',
		'clears',
		'require',
		'links',
		'connected',
		'standing',
		'wringing',
		'moaning',
		'broke',
		'querulous',
		'cry',
		'robbed',
		'helped',
		'downstairs',
		'called',
		'suspected',
		'jerked',
		'stamped',
		'convulsive',
		'frenzy',
		'report',
		'assist',
		'obeyed',
		'stumbling',
		'rubbing',
		'err',
		'underlying',
		'ejaculated',
		'clinical',
		'professor',
		'expounding',
		'class',
		'sit',
		'footprints',
		'complicate',
		'matters',
		'folk',
		'carried',
		'muttering',
		'aloud',
		'snibbed',
		'solid',
		'hinges',
		'reach',
		'rained',
		'print',
		'sill',
		'floor',
		'discs',
		'stump',
		'boot',
		'metal',
		'heel',
		'efficient',
		'ally',
		'scale',
		'shone',
		'brightly',
		'angle',
		'sixty',
		'ground',
		'foothold',
		'crevice',
		'aid',
		'stout',
		'securing',
		'hook',
		'active',
		'swarm',
		'depart',
		'draw',
		'untie',
		'shut',
		'snib',
		'originally',
		'minor',
		'noted',
		'fingering',
		'climber',
		'sailor',
		'horny',
		'discloses',
		'velocity',
		'becomes',
		'lifts',
		'breaks',
		'fresh',
		'annals',
		'crime',
		'themselves',
		'memory',
		'serves',
		'grate',
		'considered',
		'persisted',
		'apply',
		'precept',
		'shaking',
		'eliminated',
		'chimney',
		'roof',
		'extend',
		'researches',
		'seizing',
		'rafter',
		'lying',
		'beam',
		'apex',
		'shell',
		'furniture',
		'sloping',
		'leads',
		'press',
		'gentle',
		'startled',
		'surprised',
		'thickly',
		'prints',
		'defined',
		'perfectly',
		'scarce',
		'ordinary',
		'whisper',
		'horrid',
		'staggered',
		'failed',
		'foretell',
		'learned',
		'eagerly',
		'regained',
		'impatience',
		'compare',
		'results',
		'conceive',
		'tape',
		'measure',
		'measuring',
		'comparing',
		'examining',
		'inches',
		'planks',
		'beady',
		'gleaming',
		'bird',
		'swift',
		'furtive',
		'movements',
		'scent',
		'energy',
		'law',
		'exerting',
		'defence',
		'hunted',
		'loud',
		'crow',
		'delight',
		'misfortune',
		'tread',
		'creosote',
		'outline',
		'edge',
		'mess',
		'carboy',
		'cracked',
		'stuff',
		'leaked',
		'dog',
		'pack',
		'track',
		'trailed',
		'herring',
		'shire',
		'hound',
		'smell',
		'sounds',
		'accredited',
		'clamour',
		'voices',
		'audible',
		'below',
		'hall',
		'crash',
		'muscles',
		'state',
		'exceeding',
		'usual',
		'distortion',
		'writers',
		'vegetable',
		'alkaloid',
		'substance',
		'produce',
		'tetanus',
		'getting',
		'poison',
		'system',
		'driven',
		'erect',
		'gingerly',
		'glazed',
		'gummy',
		'dried',
		'blunt',
		'trimmed',
		'rounded',
		'knife',
		'auxiliary',
		'forces',
		'retreat',
		'nearer',
		'loudly',
		'portly',
		'suit',
		'strode',
		'burly',
		'plethoric',
		'swollen',
		'puffy',
		'pouches',
		'closely',
		'inspector',
		'uniform',
		'husky',
		'recollect',
		'wheezed',
		'theorist',
		'lectured',
		'jewel',
		'guidance',
		'lucky',
		'theorise',
		'dryly',
		'deny',
		'hit',
		'nail',
		'fastened',
		'flashes',
		'sergeant',
		'confession',
		'fit',
		'flaw',
		'slept',
		'disturbed',
		'weaving',
		'web',
		'net',
		'begins',
		'splinter',
		'wood',
		'inscribed',
		'instrument',
		'respect',
		'fat',
		'pompously',
		'poisonous',
		'murderous',
		'activity',
		'bulk',
		'squeezed',
		'afterwards',
		'exulting',
		'shrugging',
		'shoulders',
		'pas',
		'des',
		'sots',
		'incommodes',
		'que',
		'ceux',
		'qui',
		'ont',
		'partly',
		'discovery',
		'whoever',
		'noticed',
		'gentleman',
		'inform',
		'arrest',
		'engage',
		'harder',
		'free',
		'wearing',
		'worn',
		'sole',
		'iron',
		'band',
		'sunburned',
		'convict',
		'coupled',
		'palm',
		'sneering',
		'easily',
		'precision',
		'introduce',
		'stair',
		'occurrence',
		'lose',
		'original',
		'purpose',
		'stricken',
		'lives',
		'succession',
		'surprises',
		'nerve',
		'completely',
		'exult',
		'construct',
		'weasel',
		'rabbit',
		'queer',
		'mongrel',
		'amazing',
		'help',
		'sleeps',
		'listen',
		'sarcasms',
		'sind',
		'gewohnt',
		'das',
		'die',
		'sie',
		'nicht',
		'pithy',
		'escorted',
		'angelic',
		'borne',
		'herself',
		'support',
		'placid',
		'passion',
		'distant',
		'struggle',
		'breast',
		'effort',
		'sympathies',
		'teach',
		'brave',
		'obtrude',
		'successful',
		'honourable',
		'intimacy',
		'vulgar',
		'intervened',
		'impassable',
		'barrier',
		'interested',
		'graceful',
		'tenderly',
		'waist',
		'motherly',
		'greeted',
		'paid',
		'dependant',
		'honoured',
		'introduced',
		'begged',
		'promised',
		'faithfully',
		'progress',
		'group',
		'clinging',
		'stained',
		'barometer',
		'glimpse',
		'tranquil',
		'wilder',
		'reviewed',
		'sequence',
		'tragic',
		'baggage',
		'scene',
		'discoverer',
		'weapons',
		'endowed',
		'despair',
		'row',
		'shabby',
		'upper',
		'drunken',
		'vagabone',
		'kick',
		'kennels',
		'dogs',
		'gracious',
		'wiper',
		'bag',
		'drop',
		'argued',
		'shouted',
		'goes',
		'magical',
		'slammed',
		'unbarred',
		'lanky',
		'lean',
		'stringy',
		'neck',
		'glasses',
		'bites',
		'naughty',
		'nip',
		'stoat',
		'wicked',
		'cage',
		'fangs',
		'gives',
		'run',
		'keeps',
		'beetles',
		'guyed',
		'lane',
		'wanted',
		'animal',
		'gathered',
		'uncertain',
		'shadowy',
		'dimly',
		'glancing',
		'glimmering',
		'cranny',
		'lined',
		'solemn',
		'fowls',
		'lazily',
		'shifted',
		'slumbers',
		'ugly',
		'creature',
		'spaniel',
		'lurcher',
		'clumsy',
		'waddling',
		'gait',
		'accepted',
		'hesitation',
		'lump',
		'sugar',
		'naturalist',
		'thus',
		'alliance',
		'clock',
		'arrested',
		'accessory',
		'marched',
		'constables',
		'guarded',
		'gate',
		'allowed',
		'mentioning',
		'pockets',
		'immense',
		'display',
		'gatekeeper',
		'upstairs',
		'tied',
		'central',
		'reclined',
		'tie',
		'bit',
		'boots',
		'carry',
		'climbing',
		'dip',
		'creasote',
		'clambered',
		'footmarks',
		'noteworthy',
		'belong',
		'chief',
		'toes',
		'cramped',
		'toe',
		'divided',
		'stay',
		'strong',
		'tarry',
		'difficulty',
		'enormous',
		'crawling',
		'ridge',
		'stack',
		'chimneys',
		'reappeared',
		'vanished',
		'eaves',
		'climb',
		'feels',
		'anyhow',
		'scuffling',
		'steadily',
		'barrel',
		'easy',
		'drawing',
		'stockings',
		'loosened',
		'hurry',
		'confirms',
		'diagnosis',
		'doctors',
		'express',
		'pouch',
		'woven',
		'grasses',
		'beads',
		'strung',
		'shape',
		'spines',
		'hellish',
		'prick',
		'sooner',
		'trudge',
		'pushed',
		'fluffy',
		'separated',
		'comical',
		'cock',
		'sniffing',
		'famous',
		'vintage',
		'cord',
		'tremulous',
		'yelps',
		'tail',
		'pattered',
		'trail',
		'strained',
		'leash',
		'speed',
		'east',
		'gradually',
		'massive',
		'empty',
		'windows',
		'bare',
		'towered',
		'sad',
		'forlorn',
		'trenches',
		'pits',
		'scattered',
		'shrubs',
		'blighted',
		'harmonized',
		'tragedy',
		'boundary',
		'whining',
		'underneath',
		'screened',
		'beech',
		'bricks',
		'crevices',
		'frequently',
		'ladder',
		'smudge',
		'rain',
		'lie',
		'reflected',
		'traffic',
		'interval',
		'fears',
		'appeased',
		'hesitated',
		'swerved',
		'waddled',
		'rolling',
		'contending',
		'scents',
		'success',
		'fellows',
		'enable',
		'different',
		'ways',
		'readiest',
		'fortune',
		'culpable',
		'neglected',
		'prevented',
		'becoming',
		'gained',
		'palpable',
		'spare',
		'marvel',
		'obtain',
		'describe',
		'theatrical',
		'patent',
		'buried',
		'map',
		'named',
		'chart',
		'signed',
		'behalf',
		'brings',
		'condition',
		'dated',
		'convicts',
		'associates',
		'hypothesis',
		'covers',
		'sequel',
		'fright',
		'escaped',
		'term',
		'guards',
		'mistakes',
		'fires',
		'pistol',
		'others',
		'identical',
		'strike',
		'concise',
		'regaining',
		'consider',
		'revenge',
		'possibly',
		'butler',
		'hid',
		'learns',
		'lest',
		'runs',
		'gauntlet',
		'makes',
		'dying',
		'deterred',
		'hate',
		'enters',
		'searches',
		'private',
		'memorandum',
		'relating',
		'momento',
		'visit',
		'doubtless',
		'planned',
		'beforehand',
		'slay',
		'record',
		'bizarre',
		'conceits',
		'continue',
		'efforts',
		'household',
		'lofty',
		'takes',
		'associate',
		'gets',
		'dips',
		'whence',
		'limp',
		'damaged',
		'tendo',
		'committed',
		'disgust',
		'grudge',
		'preferred',
		'simply',
		'bound',
		'gagged',
		'halter',
		'savage',
		'instincts',
		'decipher',
		'serving',
		'oven',
		'calculated',
		'stride',
		'hairiness',
		'cloud',
		'floats',
		'pink',
		'flamingo',
		'rim',
		'sun',
		'pushes',
		'shines',
		'bet',
		'stranger',
		'ambitions',
		'strivings',
		'elemental',
		'following',
		'brook',
		'parent',
		'lake',
		'profound',
		'real',
		'greatness',
		'perception',
		'smallness',
		'argues',
		'comparison',
		'nobility',
		'food',
		'lair',
		'turns',
		'nasty',
		'shoot',
		'loaded',
		'chambers',
		'jacket',
		'roads',
		'metropolis',
		'beginning',
		'labourers',
		'dockmen',
		'astir',
		'slatternly',
		'shutters',
		'brushing',
		'emerging',
		'sleeves',
		'beards',
		'wet',
		'sauntered',
		'inimitable',
		'trotted',
		'onwards',
		'whine',
		'traversed',
		'pursued',
		'curiously',
		'zigzag',
		'escaping',
		'main',
		'edged',
		'latter',
		'advance',
		'forwards',
		'cocked',
		'canine',
		'indecision',
		'sympathy',
		'deuce',
		'growled',
		'balloon',
		'relief',
		'darted',
		'shown',
		'hotter',
		'tugged',
		'gleam',
		'nearing',
		'tavern',
		'frantic',
		'excitement',
		'enclosure',
		'sawyers',
		'raced',
		'sawdust',
		'shavings',
		'alley',
		'triumphant',
		'yelp',
		'lolling',
		'tongue',
		'blinking',
		'cask',
		'staves',
		'trolley',
		'smeared',
		'blankly',
		'laughter',
		'acted',
		'according',
		'lights',
		'lifting',
		'carted',
		'crossed',
		'seasoning',
		'blame',
		'puzzled',
		'trails',
		'leading',
		'cast',
		'circle',
		'whereas',
		'roadway',
		'tended',
		'wharf',
		'current',
		'boat',
		'punts',
		'skiffs',
		'sniffed',
		'rude',
		'placard',
		'slung',
		'printed',
		'hire',
		'steam',
		'launch',
		'pile',
		'coke',
		'jetty',
		'ominous',
		'sharper',
		'tracks',
		'management',
		'lad',
		'stoutish',
		'sponge',
		'washed',
		'finds',
		'pondered',
		'prodigy',
		'manage',
		'yesterday',
		'maybe',
		'puzzles',
		'coals',
		'barge',
		'job',
		'stayed',
		'prices',
		'odd',
		'bags',
		'outlandish',
		'talk',
		'bland',
		'chap',
		'tapped',
		'woke',
		'stones',
		'reports',
		'green',
		'trim',
		'painted',
		'streaks',
		'uneasy',
		'funnel',
		'sides',
		'boatman',
		'wherry',
		'sheets',
		'oyster',
		'colossal',
		'task',
		'touched',
		'miles',
		'exhaust',
		'injure',
		'working',
		'advertise',
		'chase',
		'push',
		'runaways',
		'landed',
		'hansom',
		'breakfast',
		'sleep',
		'cards',
		'afoot',
		'despatched',
		'resumed',
		'dirty',
		'lieutenant',
		'gang',
		'eight',
		'nine',
		'successive',
		'befogged',
		'fatigued',
		'enthusiasm',
		'antipathy',
		'murderers',
		'rightfully',
		'recovering',
		'ready',
		'devote',
		'forever',
		'selfish',
		'influenced',
		'tenfold',
		'stronger',
		'urge',
		'bath',
		'freshened',
		'coffee',
		'pointing',
		'energetic',
		'ubiquitous',
		'reporter',
		'ham',
		'eggs',
		'headed',
		'foul',
		'play',
		'actual',
		'violence',
		'gems',
		'deceased',
		'member',
		'alarm',
		'faculties',
		'gratifying',
		'result',
		'thief',
		'thieves',
		'acquainted',
		'miscreants',
		'proves',
		'haphazard',
		'burglary',
		'prompt',
		'occasions',
		'vigorous',
		'masterful',
		'supplies',
		'argument',
		'detectives',
		'closer',
		'effective',
		'grinning',
		'shave',
		'safety',
		'happen',
		'attacks',
		'ring',
		'bell',
		'wail',
		'dismay',
		'heaven',
		'irregulars',
		'pattering',
		'clatter',
		'ragged',
		'discipline',
		'despite',
		'tumultuous',
		'entry',
		'facing',
		'expectant',
		'taller',
		'older',
		'lounging',
		'funny',
		'scarecrow',
		'bob',
		'tanner',
		'tickets',
		'invaded',
		'owner',
		'boy',
		'divide',
		'banks',
		'thoroughly',
		'guinea',
		'shilling',
		'buzzed',
		'overhear',
		'spotted',
		'meanwhile',
		'await',
		'eat',
		'scraps',
		'tired',
		'idleness',
		'exhausts',
		'ours',
		'unique',
		'anyway',
		'fettered',
		'mace',
		'agility',
		'darts',
		'signs',
		'thong',
		'commonly',
		'hazarded',
		'stretched',
		'bulky',
		'shelf',
		'gazetteer',
		'authority',
		'situated',
		'north',
		'climate',
		'coral',
		'reefs',
		'sharks',
		'aborigines',
		'smallest',
		'race',
		'del',
		'average',
		'adults',
		'smaller',
		'morose',
		'capable',
		'forming',
		'hideous',
		'misshapen',
		'distorted',
		'remarkably',
		'win',
		'degree',
		'crews',
		'braining',
		'survivors',
		'clubs',
		'arrows',
		'massacres',
		'invariably',
		'concluded',
		'cannibal',
		'unaided',
		'devices',
		'affair',
		'islander',
		'regularly',
		'sofa',
		'violin',
		'melodious',
		'gift',
		'gaunt',
		'earnest',
		'fall',
		'bow',
		'floated',
		'peacefully',
		'sea',
		'dreamland',
		'refreshed',
		'aside',
		'book',
		'stirred',
		'troubled',
		'soundly',
		'wake',
		'definite',
		'provoking',
		'check',
		'outing',
		'absence',
		'twinkle',
		'pause',
		'argue',
		'atrocious',
		'sentiment',
		'curiosity',
		'dreadful',
		'parts',
		'method',
		'omissions',
		'startle',
		'amaze',
		'injured',
		'ruffian',
		'dragon',
		'earl',
		'rescue',
		'depends',
		'issue',
		'elation',
		'prospect',
		'toss',
		'behaved',
		'honourably',
		'throughout',
		'unfounded',
		'seeing',
		'note',
		'blinds',
		'sinking',
		'impressive',
		'afraid',
		'footstep',
		'talking',
		'rang',
		'stairhead',
		'cooling',
		'medicine',
		'worthy',
		'spirit',
		'chafing',
		'inaction',
		'fleck',
		'feverish',
		'cheek',
		'marching',
		'infernal',
		'consuming',
		'balked',
		'overcome',
		'disposal',
		'husband',
		'scuttled',
		'craft',
		'objections',
		'dismissed',
		'articles',
		'hostile',
		'inquest',
		'ladies',
		'dejected',
		'busied',
		'heating',
		'distilling',
		'vapours',
		'ending',
		'clinking',
		'malodorous',
		'experiment',
		'early',
		'dawn',
		'bedside',
		'scarf',
		'trying',
		'useful',
		'loath',
		'despondent',
		'telegrams',
		'allusion',
		'promises',
		'complex',
		'evidence',
		'released',
		'culprits',
		'prosecuted',
		'arrests',
		'rate',
		'whenever',
		'blunder',
		'caught',
		'agony',
		'stripes',
		'pounds',
		'doing',
		'ingenious',
		'fugitives',
		'wife',
		'imagined',
		'returning',
		'wander',
		'villainous',
		'pursuing',
		'wondered',
		'radical',
		'nimble',
		'built',
		'faulty',
		'keenest',
		'reasoner',
		'deceived',
		'error',
		'preference',
		'plainer',
		'reasons',
		'deductions',
		'trivial',
		'tending',
		'disguise',
		'incorrect',
		'equally',
		'startling',
		'peal',
		'brusque',
		'meek',
		'apologetic',
		'cigars',
		'mopping',
		'bandanna',
		'worry',
		'expressed',
		'obliged',
		'pop',
		'middle',
		'alibi',
		'climbed',
		'roofs',
		'stake',
		'jumping',
		'promising',
		'finish',
		'evident',
		'slip',
		'ascending',
		'wheezing',
		'twice',
		'aged',
		'seafaring',
		'garb',
		'bowed',
		'shaky',
		'painfully',
		'asthmatic',
		'oaken',
		'cudgel',
		'heaved',
		'lungs',
		'chin',
		'bushy',
		'brows',
		'mariner',
		'fallen',
		'acting',
		'petulant',
		'obstinacy',
		'shuffled',
		'walk',
		'returns',
		'recognised',
		'resistance',
		'stamping',
		'seize',
		'treat',
		'recompense',
		'sullenly',
		'cigar',
		'chairs',
		'sitting',
		'whiskers',
		'actor',
		'workhouse',
		'cough',
		'lighting',
		'classes',
		'publishing',
		'release',
		'prisoners',
		'fast',
		'managed',
		'telephone',
		'stanch',
		'belongs',
		'proceeding',
		'wink',
		'detail',
		'elsewhere',
		'refuse',
		'understood',
		'insist',
		'dining',
		'oysters',
		'brace',
		'grouse',
		'choice',
		'merits',
		'meal',
		'chose',
		'brilliant',
		'pottery',
		'violins',
		'humour',
		'preceding',
		'sociable',
		'relaxation',
		'faced',
		'dinner',
		'elated',
		'gaiety',
		'alluded',
		'cloth',
		'cleared',
		'port',
		'bumper',
		'prepared',
		'ordered',
		'eyed',
		'critically',
		'ropes',
		'stern',
		'rudder',
		'tend',
		'engines',
		'barges',
		'stationary',
		'overhauled',
		'steamer',
		'launches',
		'clipper',
		'land',
		'thorough',
		'plunging',
		'statesmen',
		'dissolving',
		'boys',
		'cunning',
		'finesse',
		'product',
		'education',
		'continual',
		'arrange',
		'affairs',
		'probable',
		'arranged',
		'reserved',
		'escape',
		'lodgings',
		'couple',
		'nights',
		'ship',
		'pursuit',
		'shoes',
		'repairer',
		'trifling',
		'removed',
		'shed',
		'yard',
		'liable',
		'overlooked',
		'rig',
		'inquired',
		'yards',
		'blank',
		'fifteen',
		'naught',
		'foreman',
		'liquor',
		'bellowed',
		'flush',
		'chucking',
		'shillings',
		'subsided',
		'happening',
		'stationed',
		'sentry',
		'wave',
		'neatly',
		'shrewd',
		'scout',
		'ahead',
		'suspicious',
		'snug',
		'messages',
		'series',
		'bridges',
		'span',
		'rays',
		'gilding',
		'summit',
		'twilight',
		'masts',
		'rigging',
		'string',
		'lighters',
		'shore',
		'policemen',
		'stokers',
		'granted',
		'yonder',
		'gaslight',
		'rascals',
		'immortal',
		'spark',
		'enigma',
		'calls',
		'individual',
		'puzzle',
		'aggregate',
		'certainty',
		'vary',
		'constant',
		'flutter',
		'engineer',
		'forgive',
		'unseen',
		'flying',
		'tremendous',
		'gravely',
		'burn',
		'furnaces',
		'whizzed',
		'clanked',
		'metallic',
		'steep',
		'prow',
		'waves',
		'throb',
		'living',
		'bows',
		'flickering',
		'blur',
		'swirl',
		'foam',
		'flashed',
		'steamers',
		'hailed',
		'thundered',
		'glow',
		'aquiline',
		'pound',
		'gain',
		'minutes',
		'evil',
		'tug',
		'tow',
		'blundered',
		'helm',
		'avoided',
		'collision',
		'recover',
		'starlit',
		'boilers',
		'frail',
		'vibrated',
		'rounding',
		'resolved',
		'deck',
		'mass',
		'tiller',
		'furnace',
		'stripped',
		'shovelling',
		'winding',
		'paces',
		'coursed',
		'creatures',
		'countries',
		'checkered',
		'career',
		'sport',
		'mad',
		'panting',
		'machinery',
		'crouched',
		'busy',
		'lengths',
		'boats',
		'melancholy',
		'hail',
		'clinched',
		'fists',
		'cursing',
		'poising',
		'astride',
		'thigh',
		'downwards',
		'strident',
		'cries',
		'movement',
		'huddled',
		'tangled',
		'wrapped',
		'ulster',
		'blanket',
		'sleepless',
		'deeply',
		'bestiality',
		'cruelty',
		'glowed',
		'grinned',
		'chattered',
		'fury',
		'raises',
		'quarry',
		'apart',
		'shrieking',
		'curses',
		'unhallowed',
		'dwarf',
		'gnashing',
		'plucked',
		'covering',
		'clapped',
		'pistols',
		'whirled',
		'sideways',
		'venomous',
		'menacing',
		'amid',
		'waters',
		'southern',
		'bank',
		'clearing',
		'expanse',
		'pools',
		'stagnant',
		'beds',
		'decaying',
		'vegetation',
		'thud',
		'fugitive',
		'sodden',
		'soil',
		'struggled',
		'rage',
		'kicked',
		'mud',
		'struggles',
		'bored',
		'pin',
		'sticky',
		'alongside',
		'firmly',
		'anchored',
		'haul',
		'drag',
		'fish',
		'aboard',
		'meekly',
		'commanded',
		'hauled',
		'contained',
		'cabin',
		'steamed',
		'ooze',
		'bottom',
		'bones',
		'shores',
		'hatchway',
		'shrugged',
		'sick',
		'captive',
		'network',
		'wrinkles',
		'mahogany',
		'prominence',
		'curly',
		'unpleasing',
		'aggressive',
		'handcuffed',
		'lap',
		'rigid',
		'frankly',
		'swing',
		'grieved',
		'welted',
		'devil',
		'slack',
		'undo',
		'pull',
		'flask',
		'overpower',
		'hoped',
		'supper',
		'knifing',
		'lagged',
		'acts',
		'quickly',
		'scrambled',
		'club',
		'malice',
		'bitter',
		'nigh',
		'spend',
		'breakwater',
		'digging',
		'drains',
		'merchant',
		'curse',
		'owned',
		'guilt',
		'slavery',
		'party',
		'overhaul',
		'ends',
		'fastest',
		'swears',
		'flier',
		'vessel',
		'condemning',
		'amusing',
		'airs',
		'strength',
		'capture',
		'played',
		'speech',
		'pity',
		'inventory',
		'shortly',
		'warn',
		'bluff',
		'genial',
		'obliging',
		'diaphanous',
		'material',
		'scarlet',
		'shaded',
		'basket',
		'playing',
		'tinting',
		'sparkle',
		'coils',
		'luxuriant',
		'pose',
		'absorbing',
		'dreamed',
		'speaking',
		'jovially',
		'coolly',
		'thousand',
		'annuity',
		'richer',
		'overacting',
		'detected',
		'hollow',
		'owe',
		'taxed',
		'narrated',
		'briefly',
		'recital',
		'dart',
		'narrowly',
		'missed',
		'hastened',
		'pour',
		'peril',
		'gloomy',
		'brighter',
		'eagerness',
		'ungracious',
		'prize',
		'raise',
		'borrow',
		'poker',
		'hasp',
		'wrought',
		'image',
		'lever',
		'lid',
		'gazing',
		'price',
		'shred',
		'crumb',
		'jewelry',
		'calmly',
		'realised',
		'weighed',
		'disloyal',
		'realise',
		'withdraw',
		'truly',
		'loved',
		'whispered',
		'patient',
		'rejoined',
		'clouded',
		'gloomily',
		'tenner',
		'rewarded',
		'forecast',
		'prisoner',
		'changed',
		'plans',
		'lounged',
		'listless',
		'stolidly',
		'exhibited',
		'angrily',
		'exultantly',
		'loot',
		'darned',
		'kith',
		'kin',
		'rupees',
		'deceiving',
		'sternly',
		'easier',
		'sidelong',
		'hunt',
		'grieving',
		'ups',
		'downs',
		'spilled',
		'milk',
		'thwarting',
		'trial',
		'snarled',
		'earned',
		'swamp',
		'chained',
		'filthy',
		'bitten',
		'mosquitoes',
		'racked',
		'ague',
		'bullied',
		'enjoy',
		'score',
		'cell',
		'palace',
		'mask',
		'stoicism',
		'whirl',
		'blazed',
		'handcuffs',
		'groundless',
		'thank',
		'bracelets',
		'wrists',
		'dry',
		'steady',
		'farmers',
		'respected',
		'rover',
		'eighteen',
		'girl',
		'joining',
		'starting',
		'destined',
		'soldiering',
		'fool',
		'swimming',
		'company',
		'swimmers',
		'crocodile',
		'nipped',
		'drowned',
		'paddled',
		'hospital',
		'timber',
		'strapped',
		'invalided',
		'unfitted',
		'occupation',
		'useless',
		'cripple',
		'twentieth',
		'blessing',
		'overseer',
		'coolies',
		'accident',
		'colonel',
		'strongly',
		'mostly',
		'horseback',
		'grip',
		'saddle',
		'ride',
		'plantation',
		'idlers',
		'quarters',
		'content',
		'remainder',
		'shanty',
		'warning',
		'mutiny',
		'month',
		'peaceful',
		'devils',
		'hell',
		'reading',
		'border',
		'alight',
		'burning',
		'bungalows',
		'companies',
		'estate',
		'wives',
		'nearest',
		'obstinate',
		'veranda',
		'cheroots',
		'managing',
		'riding',
		'nullah',
		'rode',
		'ribbons',
		'eaten',
		'jackals',
		'reined',
		'curling',
		'bungalow',
		'flames',
		'meddled',
		'hundreds',
		'fiends',
		'coats',
		'backs',
		'dancing',
		'bullets',
		'sang',
		'bees',
		'collect',
		'bands',
		'guns',
		'fight',
		'millions',
		'cruellest',
		'gunners',
		'taught',
		'handling',
		'blowing',
		'battery',
		'artillery',
		'volunteer',
		'corps',
		'clerks',
		'merchants',
		'powder',
		'worst',
		'south',
		'compass',
		'torture',
		'outrage',
		'swarming',
		'fanatics',
		'sorts',
		'handful',
		'leader',
		'fort',
		'queerest',
		'rum',
		'acres',
		'garrison',
		'stores',
		'nobody',
		'scorpions',
		'centipedes',
		'deserted',
		'twisting',
		'torches',
		'exploring',
		'washes',
		'protects',
		'angles',
		'gates',
		'organise',
		'natives',
		'selected',
		'isolated',
		'southwest',
		'troopers',
		'instructed',
		'fire',
		'arrive',
		'attack',
		'raw',
		'recruit',
		'chaps',
		'jabber',
		'lingo',
		'gateway',
		'beating',
		'drums',
		'tomtoms',
		'yells',
		'howls',
		'drunk',
		'opium',
		'bang',
		'remind',
		'posts',
		'weariness',
		'match',
		'snatched',
		'firelock',
		'levelled',
		'swore',
		'plunge',
		'league',
		'assault',
		'intention',
		'scream',
		'braced',
		'noise',
		'rebel',
		'fiercer',
		'silenced',
		'hesitate',
		'oath',
		'ditch',
		'brothers',
		'truck',
		'countrymen',
		'swear',
		'threefold',
		'honour',
		'tale',
		'stands',
		'binding',
		'sworn',
		'gods',
		'temples',
		'rajah',
		'northern',
		'provinces',
		'wealth',
		'lands',
		'hoards',
		'gold',
		'troubles',
		'lion',
		'overthrow',
		'vaults',
		'precious',
		'choicest',
		'trusty',
		'guise',
		'won',
		'conquered',
		'saved',
		'hoard',
		'borders',
		'due',
		'salt',
		'pretended',
		'travels',
		'lonely',
		'sacred',
		'meeting',
		'stare',
		'moidores',
		'commandant',
		'government',
		'rupee',
		'coffers',
		'chiefs',
		'handing',
		'devised',
		'falling',
		'season',
		'drifting',
		'moat',
		'challenge',
		'uncover',
		'stopping',
		'advancing',
		'scramble',
		'splash',
		'mire',
		'challenged',
		'subdued',
		'uncovered',
		'flood',
		'beard',
		'swept',
		'cummerbund',
		'shawl',
		'quiver',
		'twitched',
		'mouse',
		'ventures',
		'chills',
		'killing',
		'flint',
		'chirrup',
		'travelled',
		'seek',
		'shelter',
		'beaten',
		'abused',
		'blessed',
		'governor',
		'compassed',
		'measured',
		'tramp',
		'sounding',
		'scuffle',
		'blows',
		'rush',
		'smear',
		'bounding',
		'flashing',
		'gaining',
		'softened',
		'stagger',
		'uttered',
		'moan',
		'muscle',
		'telling',
		'favour',
		'manacled',
		'brewed',
		'conceived',
		'flippant',
		'punishment',
		'store',
		'defiance',
		'proceeded',
		'refused',
		'throats',
		'pains',
		'lenient',
		'crumbling',
		'attacked',
		'silken',
		'carved',
		'gleamed',
		'blinding',
		'feasted',
		'list',
		'diamonds',
		'including',
		'largest',
		'emeralds',
		'rubies',
		'carbuncles',
		'sapphires',
		'agates',
		'quantity',
		'beryls',
		'onyxes',
		'turquoises',
		'familiar',
		'coronet',
		'counted',
		'treasures',
		'solemnly',
		'renewed',
		'agreed',
		'dividing',
		'privacy',
		'frontier',
		'settling',
		'safely',
		'shares',
		'plunder',
		'shattered',
		'spy',
		'refuge',
		'admission',
		'guides',
		'fourth',
		'murdered',
		'deposed',
		'penal',
		'servitude',
		'condemned',
		'commuted',
		'cuff',
		'rice',
		'gorgeous',
		'stubborn',
		'bided',
		'settlement',
		'privileged',
		'hut',
		'slopes',
		'clearings',
		'infested',
		'ditching',
		'drugs',
		'smattering',
		'lookout',
		'seas',
		'terribly',
		'sporting',
		'surgery',
		'lonesome',
		'fond',
		'crafty',
		'nice',
		'sly',
		'soldiers',
		'civilians',
		'unfair',
		'poorer',
		'hardest',
		'big',
		'sums',
		'deals',
		'thunder',
		'raving',
		'losses',
		'saying',
		'ruined',
		'slapping',
		'facer',
		'strolling',
		'beach',
		'cheroot',
		'shortened',
		'gasped',
		'outlawed',
		'rash',
		'repent',
		'changes',
		'identify',
		'stock',
		'twitch',
		'rings',
		'concern',
		'disposing',
		'agree',
		'bargain',
		'freedom',
		'theirs',
		'bar',
		'voyage',
		'provisions',
		'yachts',
		'yawls',
		'coast',
		'flinch',
		'monthly',
		'inquire',
		'growing',
		'colder',
		'consent',
		'comrades',
		'provide',
		'charts',
		'yacht',
		'duties',
		'oaths',
		'utter',
		'impatient',
		'stowed',
		'chokey',
		'villain',
		'passengers',
		'uncle',
		'stoop',
		'scoundrel',
		'carrying',
		'conditions',
		'sold',
		'vengeance',
		'nursed',
		'cared',
		'gallows',
		'slaying',
		'fever',
		'woods',
		'snake',
		'fonder',
		'roomy',
		'canoe',
		'gourds',
		'lot',
		'yams',
		'potatoes',
		'mate',
		'chanced',
		'vile',
		'insulting',
		'injuring',
		'vowed',
		'debt',
		'island',
		'carbine',
		'brains',
		'weapon',
		'unstrapped',
		'hops',
		'skull',
		'split',
		'earthly',
		'bamboo',
		'spear',
		'sail',
		'trusting',
		'eleventh',
		'trader',
		'cargo',
		'pilgrims',
		'chum',
		'drifted',
		'dream',
		'someone',
		'besides',
		'clutches',
		'bethought',
		'met',
		'token',
		'befooled',
		'exhibiting',
		'fairs',
		'meat',
		'dance',
		'hatful',
		'pennies',
		'hunting',
		'cat',
		'strutting',
		'peacock',
		'imp',
		'slid',
		'waterman',
		'screw',
		'secrets',
		'badly',
		'innocent',
		'fitting',
		'affably',
		'humoured',
		'waits',
		'inspectors',
		'wary',
		'drama',
		'studying',
		'groan',
		'hurt',
		'charming',
		'decided',
		'witness',
		'preserved',
		'opposed',
		'marry',
		'bias',
		'survive',
		'ordeal',
		'rag',
		'laziness',
		'alternate',
		'splendid',
		'vigour',
		'makings',
		'loafer',
		'spry',
		'dass',
		'nur',
		'aus',
		'schuf',
		'zum',
		'war',
		'und',
		'der',
		'surmised',
		'undivided',
		'file',
		'various',
		'formats',
		'editions',
		'replace',
		'previous',
		'renamed',
		'protected',
		'copyright',
		'owns',
		'distribute',
		'permission',
		'paying',
		'royalties',
		'rules',
		'license',
		'copying',
		'electronic',
		'protect',
		'concept',
		'trademark',
		'receive',
		'specific',
		'copies',
		'complying',
		'creation',
		'derivative',
		'modified',
		'commercial',
		'mission',
		'promoting',
		'using',
		'comply',
		'available',
		'indicate',
		'abide',
		'cease',
		'destroy',
		'fee',
		'obtaining',
		'access',
		'refund',
		'entity',
		'paragraph',
		'preserve',
		'domain',
		'located',
		'performing',
		'displaying',
		'creating',
		'based',
		'sharing',
		'compliance',
		'format',
		'attached',
		'laws',
		'govern',
		'addition',
		'concerning',
		'status',
		'immediate',
		'accessed',
		'displayed',
		'performed',
		'viewed',
		'copied',
		'ebook',
		'derived',
		'texts',
		'indicating',
		'posted',
		'fees',
		'charges',
		'providing',
		'appearing',
		'paragraphs',
		'holder',
		'imposed',
		'linked',
		'unlink',
		'detach',
		'remove',
		'perform',
		'convert',
		'binary',
		'compressed',
		'processing',
		'hypertext',
		'version',
		'site',
		'expense',
		'user',
		'exporting',
		'include',
		'specified',
		'viewing',
		'reasonable',
		'royalty',
		'gross',
		'profits',
		'derive',
		'calculate',
		'applicable',
		'taxes',
		'owed',
		'donate',
		'payments',
		'legally',
		'required',
		'periodic',
		'donations',
		'notifies',
		'receipt',
		'physical',
		'medium',
		'accordance',
		'defect',
		'reported',
		'volunteers',
		'employees',
		'expend',
		'transcribe',
		'proofread',
		'stored',
		'incomplete',
		'inaccurate',
		'corrupt',
		'errors',
		'defective',
		'disk',
		'computer',
		'virus',
		'codes',
		'damage',
		'equipment',
		'disclaim',
		'liability',
		'damages',
		'costs',
		'expenses',
		'legal',
		'elect',
		'lieu',
		'fix',
		'states',
		'implied',
		'warranties',
		'exclusion',
		'limitation',
		'types',
		'disclaimer',
		'violates',
		'maximum',
		'permitted',
		'invalidity',
		'provision',
		'void',
		'remaining',
		'indemnify',
		'agent',
		'employee',
		'production',
		'promotion',
		'arise',
		'directly',
		'indirectly',
		'occur',
		'alteration',
		'additions',
		'deletions',
		'synonymous',
		'readable',
		'widest',
		'computers',
		'obsolete',
		'exists',
		'walks',
		'financial',
		'critical',
		'goals',
		'ensuring',
		'page',
		'non',
		'profit',
		'organized',
		'exempt',
		'federal',
		'deductible',
		'principal',
		'office',
		'mailing',
		'locations',
		'increasing',
		'licensed',
		'machine',
		'accessible',
		'array',
		'outdated',
		'regulating',
		'charities',
		'charitable',
		'paperwork',
		'solicit',
		'determine',
		'accepting',
		'donors',
		'approach',
		'offers',
		'gratefully',
		'statements',
		'pages',
		'donation',
		'addresses',
		'checks',
		'originator',
		'library',
		'shared',
		'edition',
		'facility',
		'includes',
		'subscribe',
		'email',
		'newsletter',
	]
}
